`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Dennis Porras, David Gómez and Kelvin Alfaro
// 
// Create Date:    14:51:08 09/06/2017 
// Design Name: 	Modulo de Parametros
// Module Name:    Parameters 
// Project Name: Train Controller
// Target Devices: FPGA
// Tool versions: 1.0
// Description: Modulo para la verificacion de parámetros
//
// Dependencies: 
//
// Revision: 1
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Parameters(
    input A,
    input B,
    input C,
    input D,
    output T
    );


endmodule
